module LED(led);
	output led;
	
	assign led=4'b1010;
	


endmodule